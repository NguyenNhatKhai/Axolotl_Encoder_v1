////////////////////////////////////////////////////////////////////////////////////////////////////

`include "encoder.vh"

////////////////////////////////////////////////////////////////////////////////////////////////////

module enc_buffer (
    input clk,
    input rst_n,
    input con_stall,
    input [ENC_SYM_NUM - 1 : 0][EGF_ORDER - 1 : 0] enc_data,
    output logic [2 * ENC_SYM_NUM - 1 : 0][EGF_ORDER - 1 : 0] buf_data
);

////////////////////////////////////////////////////////////////////////////////////////////////////

    always_ff @(posedge clk) begin
        if (!rst_n) begin
            buf_data <= '0;
        end else if (!con_stall) begin
            buf_data[2 * ENC_SYM_NUM - 1 : ENC_SYM_NUM] <= buf_data[ENC_SYM_NUM - 1 : 0];
            buf_data[ENC_SYM_NUM - 1 : 0] <= enc_data;
        end
    end

endmodule

////////////////////////////////////////////////////////////////////////////////////////////////////